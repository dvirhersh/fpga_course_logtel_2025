--------------------------------------------------------------------------------
-- File       : demo_tb.vhd
-- Author     : AMD Inc.
--------------------------------------------------------------------------------
-- (c) Copyright 2002-2008 Advanced Micro Devices, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 
-- 
-- 
--------------------------------------------------------------------------------
--
-- Description: This test fixture will exercise the ports of the
-- Ethernet 1000BASE-X PCS/PMA core's example design to perform the
-- following operations:
--
------------------
--  Transmitter
------------------
--  Four frames are generated by the Tx Stimulus and pushed into the
--  GMII transmitter.
--
--  The PHY side transmitter interface data is captured, 8B10B decoded
--  and the Tx Monitor checks that the captured data matches that
--  injected.
--
------------------
--  Receiver
------------------
--  Four frames are generated by the Rx Stimulus, 8B10B encoded and
--  pushed into the PHY side receiver interface.
--
--  The GMII side receiver interface data is captured and the
--  Rx Monitor checks that the captured data matches that injected.


------------------------------------------------------------------------
--                    Demonstration Testbench                          |
--                                                                     |
--                                                                     |
--                  --------------------------                         |
--                  |     Example Design     |                         |
--                  |         (DUT)          |                         |
--                  |                        |                         |
--                  |                        |                         |
--                  |                        |                         |
--   Tx             |                        |  8B10B decode, Tx       |
--   Generate   ------->                  -------->           Monitor  |
--   Frames         |                        |                Frames   |
--                  |                        |                         |
--                  |GMII                PHY |                         |
--                  | I/F                I/F |                         |
--                  |                        |                         |
--                  |                        |                         |
--    Rx            |                        |  8B10B encode, Rx       |
--    Monitor  <--------                  <--------           Generate |
--    Frames        |                        |                Frames   |
--                  |                        |                         |
--                  --------------------------                         |
--                                                                     |
--                                                                     |
------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;



--------------------------------------------------------------------------------
-- This entity is the ethernet frame stimulus testbench
--------------------------------------------------------------------------------

entity stimulus_tb is
    generic (
      INSTANCE_NUMBER          : integer := 0
    );
    port (

      -- Physical Interface (TBI)
      ---------------------------
      gtx_clk                 : out std_logic;
      pma_tx_clk              : in  std_logic;
      tx_code_group           : in  std_logic_vector(9 downto 0);
      rx_code_group           : out std_logic_vector(9 downto 0);
      pma_rx_clk0             : out std_logic;
      pma_rx_clk1             : out std_logic;

      -- GMII Interface
      -----------------
      gmii_tx_clk             : out std_logic;
      gmii_rx_clk             : in std_logic;
      gmii_txd                : out std_logic_vector(7 downto 0);
      gmii_tx_en              : out std_logic;
      gmii_tx_er              : out std_logic;
      gmii_rxd                : in std_logic_vector(7 downto 0);
      gmii_rx_dv              : in std_logic;
      gmii_rx_er              : in std_logic;

      -- Test bench speed selection
      -----------------------------
      speed_is_10_100         : in std_logic;
      speed_is_100            : in std_logic;

      -- Test Bench Semaphores
      ------------------------
      configuration_finished  : in  boolean;
      tx_monitor_finished     : out boolean;
      rx_monitor_finished     : out boolean
      );
end stimulus_tb;



architecture behav of stimulus_tb is


-- Unit Interval for Gigabit Ethernet
  constant UI    : time := 800 ps;
    


  ------------------------------------------------------------------------------
  -- Procedure to perform 8B10B decoding
  ------------------------------------------------------------------------------

  -- Decode the 8B10B code. No disparity verification is performed, just
  -- a simple table lookup.
  procedure decode_8b10b (
    constant d10  : in  std_logic_vector(0 to 9);
    variable q8   : out std_logic_vector(7 downto 0);
    variable is_k : out boolean) is
    variable k28 : boolean;
    variable d10_rev : std_logic_vector(9 downto 0);
  begin
    -- reverse the 10B codeword
    for i in 0 to 9 loop
      d10_rev(i) := d10(i);
    end loop;  -- i
    -- do the 6B5B decode
    case d10_rev(5 downto 0) is
      when "000110" =>
        q8(4 downto 0) := "00000";   --D.0
      when "111001" =>
        q8(4 downto 0) := "00000";   --D.0
      when "010001" =>
        q8(4 downto 0) := "00001";   --D.1
      when "101110" =>
        q8(4 downto 0) := "00001";   --D.1
      when "010010" =>
        q8(4 downto 0) := "00010";   --D.2
      when "101101" =>
        q8(4 downto 0) := "00010";   --D.2
      when "100011" =>
        q8(4 downto 0) := "00011";   --D.3
      when "010100" =>
        q8(4 downto 0) := "00100";   --D.4
      when "101011" =>
        q8(4 downto 0) := "00100";   --D.4
      when "100101" =>
        q8(4 downto 0) := "00101";   --D.5
      when "100110" =>
        q8(4 downto 0) := "00110";   --D.6
      when "000111" =>
        q8(4 downto 0) := "00111";   --D.7
      when "111000" =>
        q8(4 downto 0) := "00111";   --D.7
      when "011000" =>
        q8(4 downto 0) := "01000";   --D.8
      when "100111" =>
        q8(4 downto 0) := "01000";   --D.8
      when "101001" =>
        q8(4 downto 0) := "01001";   --D.9
      when "101010" =>
        q8(4 downto 0) := "01010";   --D.10
      when "001011" =>
        q8(4 downto 0) := "01011";   --D.11
      when "101100" =>
        q8(4 downto 0) := "01100";   --D.12
      when "001101" =>
        q8(4 downto 0) := "01101";   --D.13
      when "001110" =>
        q8(4 downto 0) := "01110";   --D.14
      when "000101" =>
        q8(4 downto 0) := "01111";   --D.15
      when "111010" =>
        q8(4 downto 0) := "01111";   --D.15
      when "110110" =>
        q8(4 downto 0) := "10000";   --D.16
      when "001001" =>
        q8(4 downto 0) := "10000";   --D.16
      when "110001" =>
        q8(4 downto 0) := "10001";   --D.17
      when "110010" =>
        q8(4 downto 0) := "10010";   --D.18
      when "010011" =>
        q8(4 downto 0) := "10011";   --D.19
      when "110100" =>
        q8(4 downto 0) := "10100";   --D.20
      when "010101" =>
        q8(4 downto 0) := "10101";   --D.21
      when "010110" =>
        q8(4 downto 0) := "10110";   --D.22
      when "010111" =>
        q8(4 downto 0) := "10111";   --D/K.23
      when "101000" =>
        q8(4 downto 0) := "10111";   --D/K.23
      when "001100" =>
        q8(4 downto 0) := "11000";   --D.24
      when "110011" =>
        q8(4 downto 0) := "11000";   --D.24
      when "011001" =>
        q8(4 downto 0) := "11001";   --D.25
      when "011010" =>
        q8(4 downto 0) := "11010";   --D.26
      when "011011" =>
        q8(4 downto 0) := "11011";   --D/K.27
      when "100100" =>
        q8(4 downto 0) := "11011";   --D/K.27
      when "011100" =>
        q8(4 downto 0) := "11100";   --D.28
      when "111100" =>
        q8(4 downto 0) := "11100";   --K.28
      when "000011" =>
        q8(4 downto 0) := "11100";   --K.28
      when "011101" =>
        q8(4 downto 0) := "11101";   --D/K.29
      when "100010" =>
        q8(4 downto 0) := "11101";   --D/K.29
      when "011110" =>
        q8(4 downto 0) := "11110";   --D.30
      when "100001" =>
        q8(4 downto 0) := "11110";   --D.30
      when "110101" =>
        q8(4 downto 0) := "11111";   --D.31
      when "001010" =>
        q8(4 downto 0) := "11111";   --D.31

      when others   =>
        q8(4 downto 0) := "11110";  --CODE VIOLATION - return /E/
    end case;

    k28 := not((d10(2) OR d10(3) OR d10(4) OR d10(5)
                OR NOT(d10(8) XOR d10(9)))) = '1';

    -- do the 4B3B decode
    case d10_rev(9 downto 6) is
      when "0010" =>
        q8(7 downto 5) := "000";       --D/K.x.0
      when "1101" =>
        q8(7 downto 5) := "000";       --D/K.x.0
      when "1001" =>
        if not k28 then
          q8(7 downto 5) := "001";     --D/K.x.1
        else
          q8(7 downto 5) := "110";     --K28.6
        end if;
      when "0110" =>
        if k28 then
          q8(7 downto 5) := "001";     --K.28.1
        else
          q8(7 downto 5) := "110";     --D/K.x.6
        end if;
      when "1010" =>
        if not k28 then
          q8(7 downto 5) := "010";     --D/K.x.2
        else
          q8(7 downto 5) := "101";     --K28.5
        end if;
      when "0101" =>
        if k28 then
          q8(7 downto 5) := "010";     --K28.2
        else
          q8(7 downto 5) := "101";     --D/K.x.5
        end if;
      when "0011" =>
        q8(7 downto 5) := "011";       --D/K.x.3
      when "1100" =>
        q8(7 downto 5) := "011";       --D/K.x.3
      when "0100" =>
        q8(7 downto 5) := "100";       --D/K.x.4
      when "1011" =>
        q8(7 downto 5) := "100";       --D/K.x.4
      when "0111" =>
        q8(7 downto 5) := "111";       --D.x.7
      when "1000" =>
        q8(7 downto 5) := "111";       --D.x.7
      when "1110" =>
        q8(7 downto 5) := "111";       --D/K.x.7
      when "0001" =>
        q8(7 downto 5) := "111";       --D/K.x.7

      when others =>
        q8(7 downto 5) := "111";   --CODE VIOLATION - return /E/
    end case;

    is_k := ((d10(2) and d10(3) and d10(4) and d10(5))
            or not (d10(2) or d10(3) or d10(4) or d10(5))
            or ((d10(4) xor d10(5))
              and ((d10(5) and d10(7) and d10(8) and d10(9))
                or not(d10(5) or d10(7) or d10(8) or d10(9))))) = '1' ;
  end decode_8b10b;



  ------------------------------------------------------------------------------
  -- Procedure to perform comma detection
  ------------------------------------------------------------------------------

  function is_comma (
    constant codegroup : in std_logic_vector(0 to 9))
    return boolean is
  begin  -- is_comma
    case codegroup(0 to 6) is
      when "0011111" =>
        return true;
      when "1100000" =>
        return true;
      when others =>
        return false;
    end case;
  end is_comma;


  ------------------------------------------------------------------------------
  -- Procedure to perform 8B10B encoding
  ------------------------------------------------------------------------------

  procedure encode_8b10b (
    constant d8                : in  std_logic_vector(7 downto 0);
    constant is_k              : in  boolean;
    variable q10               : out std_logic_vector(0 to 9);
    constant disparity_pos_in  : in  boolean;
    variable disparity_pos_out : out boolean) is
    variable b6                       : std_logic_vector(5 downto 0);
    variable b4                       : std_logic_vector(3 downto 0);
    variable k28, pdes6, a7, l13, l31 : boolean;
    variable a, b, c, d, e            : boolean;
  begin  -- encode_8b10b
    -- precalculate some common terms
    a := d8(0) = '1';
    b := d8(1) = '1';
    c := d8(2) = '1';
    d := d8(3) = '1';
    e := d8(4) = '1';

    k28 := is_k and d8(4 downto 0) = "11100";
    l13 := (((a xor b) and not (c or d))
            or ((c xor d) and not(a or b)));

    l31 := (((a xor b) and (c and d))
             or
             ((c xor d) and (a and b)));

    a7 := is_k or ((l31 and d and not e and disparity_pos_in)
                   or (l13 and not d and e and not disparity_pos_in));

    -- Do the 5B/6B conversion (calculate the 6b symbol)
    if k28 then                         --K.28
      if not disparity_pos_in then
        b6 := "111100";
      else
        b6 := "000011";
      end if;
    else
      case d8(4 downto 0) is
        when "00000" =>                 --D.0
          if disparity_pos_in then
            b6 := "000110";
          else
            b6 := "111001";
          end if;
        when "00001" =>                 --D.1
          if disparity_pos_in then
            b6 := "010001";
          else
            b6 := "101110";
          end if;
        when "00010" =>                 --D.2
          if disparity_pos_in then
            b6 := "010010";
          else
            b6 := "101101";
          end if;
        when "00011" =>
          b6 := "100011";               --D.3
        when "00100" =>                 --D.4
          if disparity_pos_in then
            b6 := "010100";
          else
            b6 := "101011";
          end if;
        when "00101" =>
          b6 := "100101";               --D.5
        when "00110" =>
          b6 := "100110";               --D.6
        when "00111" =>                 --D.7
          if not disparity_pos_in then
            b6 := "000111";
          else
            b6 := "111000";
          end if;
        when "01000" =>                 --D.8
          if disparity_pos_in then
            b6 := "011000";
          else
            b6 := "100111";
          end if;
        when "01001" =>
          b6 := "101001";               --D.9
        when "01010" =>
          b6 := "101010";               --D.10
        when "01011" =>
          b6 := "001011";               --D.11
        when "01100" =>
          b6 := "101100";               --D.12
        when "01101" =>
          b6 := "001101";               --D.13
        when "01110" =>
          b6 := "001110";               --D.14
        when "01111" =>                 --D.15
          if disparity_pos_in then
            b6 := "000101";
          else
            b6 := "111010";
          end if;
        when "10000" =>                 --D.16
          if not disparity_pos_in then
            b6 := "110110";
          else
            b6 := "001001";
          end if;
        when "10001" =>
          b6 := "110001";               --D.17
        when "10010" =>
          b6 := "110010";               --D.18
        when "10011" =>
          b6 := "010011";               --D.19
        when "10100" =>
          b6 := "110100";               --D.20
        when "10101" =>
          b6 := "010101";               --D.21
        when "10110" =>
          b6 := "010110";               --D.22
        when "10111" =>                 --D/K.23
          if not disparity_pos_in then
            b6 := "010111";
          else
            b6 := "101000";
          end if;
        when "11000" =>                 --D.24
          if disparity_pos_in then
            b6 := "001100";
          else
            b6 := "110011";
          end if;
        when "11001" =>
          b6 := "011001";               --D.25
        when "11010" =>
          b6 := "011010";               --D.26
        when "11011" =>                 --D/K.27
          if not disparity_pos_in then
            b6 := "011011";
          else
            b6 := "100100";
          end if;
        when "11100" =>
          b6 := "011100";               --D.28
        when "11101" =>                 --D/K.29
          if not disparity_pos_in then
            b6 := "011101";
          else
            b6 := "100010";
          end if;
        when "11110" =>                 --D/K.30
          if not disparity_pos_in then
            b6 := "011110";
          else
            b6 := "100001";
          end if;
        when "11111" =>                 --D.31
          if not disparity_pos_in then
            b6 := "110101";
          else
            b6 := "001010";
          end if;
        when others =>
          b6 := "XXXXXX";
      end case;
    end if;

    -- reverse the bits
    for i in 0 to 5 loop
      q10(i) := b6(i);
    end loop;  -- i

    -- calculate the running disparity after the 5B6B block encode
    if k28 then
      pdes6 := not disparity_pos_in;
    else
      case d8(4 downto 0) is
        when "00000" => pdes6 := not disparity_pos_in;
        when "00001" => pdes6 := not disparity_pos_in;
        when "00010" => pdes6 := not disparity_pos_in;
        when "00011" => pdes6 := disparity_pos_in;
        when "00100" => pdes6 := not disparity_pos_in;
        when "00101" => pdes6 := disparity_pos_in;
        when "00110" => pdes6 := disparity_pos_in;
        when "00111" => pdes6 := disparity_pos_in;

        when "01000" => pdes6 := not disparity_pos_in;
        when "01001" => pdes6 := disparity_pos_in;
        when "01010" => pdes6 := disparity_pos_in;
        when "01011" => pdes6 := disparity_pos_in;
        when "01100" => pdes6 := disparity_pos_in;
        when "01101" => pdes6 := disparity_pos_in;
        when "01110" => pdes6 := disparity_pos_in;
        when "01111" => pdes6 := not disparity_pos_in;

        when "10000" => pdes6 := not disparity_pos_in;
        when "10001" => pdes6 := disparity_pos_in;
        when "10010" => pdes6 := disparity_pos_in;
        when "10011" => pdes6 := disparity_pos_in;
        when "10100" => pdes6 := disparity_pos_in;
        when "10101" => pdes6 := disparity_pos_in;
        when "10110" => pdes6 := disparity_pos_in;
        when "10111" => pdes6 := not disparity_pos_in;

        when "11000" => pdes6 := not disparity_pos_in;
        when "11001" => pdes6 := disparity_pos_in;
        when "11010" => pdes6 := disparity_pos_in;
        when "11011" => pdes6 := not disparity_pos_in;
        when "11100" => pdes6 := disparity_pos_in;
        when "11101" => pdes6 := not disparity_pos_in;
        when "11110" => pdes6 := not disparity_pos_in;
        when "11111" => pdes6 := not disparity_pos_in;
        when others  => pdes6 := disparity_pos_in;
      end case;
    end if;

    case d8(7 downto 5) is
      when "000" =>                     --D/K.x.0
        if pdes6 then
          b4 := "0010";
        else
          b4 := "1101";
        end if;
      when "001" =>                     --D/K.x.1
        if k28 and not pdes6 then
          b4 := "0110";
        else
          b4 := "1001";
        end if;
      when "010" =>                     --D/K.x.2
        if k28 and not pdes6 then
          b4 := "0101";
        else
          b4 := "1010";
        end if;
      when "011" =>                     --D/K.x.3
        if not pdes6 then
          b4 := "0011";
        else
          b4 := "1100";
        end if;
      when "100" =>                     --D/K.x.4
        if pdes6 then
          b4 := "0100";
        else
          b4 := "1011";
        end if;
      when "101" =>                     --D/K.x.5
        if k28 and not pdes6 then
          b4 := "1010";
        else
          b4 := "0101";
        end if;
      when "110" =>                     --D/K.x.6
        if k28 and not pdes6 then
          b4 := "1001";
        else
          b4 := "0110";
        end if;
      when "111" =>                     --D.x.P7
        if not a7 then
          if not pdes6 then
            b4 := "0111";
          else
            b4 := "1000";
          end if;
        else                            --D/K.y.A7
          if not pdes6 then
            b4 := "1110";
          else
            b4 := "0001";
          end if;
        end if;
      when others =>
        b4 := "XXXX";
    end case;

    -- Reverse the bits
    for i in 0 to 3 loop
      q10(i+6) := b4(i);
    end loop;  -- i

    -- Calculate the running disparity after the 4B group
    case d8(7 downto 5) is
      when "000"  =>
        disparity_pos_out := not pdes6;
      when "001"  =>
        disparity_pos_out := pdes6;
      when "010"  =>
        disparity_pos_out := pdes6;
      when "011"  =>
        disparity_pos_out := pdes6;
      when "100"  =>
        disparity_pos_out := not pdes6;
      when "101"  =>
        disparity_pos_out := pdes6;
      when "110"  =>
        disparity_pos_out := pdes6;
      when "111"  =>
        disparity_pos_out := not pdes6;
      when others =>
        disparity_pos_out := pdes6;
    end case;

  end encode_8b10b;



  ------------------------------------------------------------------------------
  -- types to support frame data
  ------------------------------------------------------------------------------
  -- gmii_txd, gmii_tx_en and gmii_tx_er record
  type data_typ is record
                       data  : bit_vector(7 downto 0);  -- data
                       valid : bit;                     -- data valid
                       error : bit;                     -- data error
                     end record;
  type frame_of_data_typ is array (natural range <>) of data_typ;

  -- Tx Data, Data_valid and underrun record
  type frame_typ is record
                      columns  : frame_of_data_typ(0 to 73);
                    end record;
  type frame_typ_ary is array (natural range <>) of frame_typ;



  ------------------------------------------------------------------------------
  -- Stimulus - Frame data
  ------------------------------------------------------------------------------
  -- The following constant holds the stimulus for the testbench. It is
  -- an ordered array of frames, with frame 0 the first to be injected
  -- into the core by the testbench.
  --
  -- This stimulus is used for both transmitter and receiver paths.
  ------------------------------------------------------------------------------
  constant frame_data : frame_typ_ary := (
    0          => (                     -- Frame 0
      columns  => (
        0      => ( data => X"55", valid => '1', error => '0'), -- Preamble
        1      => ( data => X"55", valid => '1', error => '0'),
        2      => ( data => X"55", valid => '1', error => '0'),
        3      => ( data => X"55", valid => '1', error => '0'),
        4      => ( data => X"55", valid => '1', error => '0'),
        5      => ( data => X"55", valid => '1', error => '0'),
        6      => ( data => X"55", valid => '1', error => '0'),
        7      => ( data => X"D5", valid => '1', error => '0'), -- SFD
        8      => ( data => X"DA", valid => '1', error => '0'), -- Destination Address (DA)
        9      => ( data => X"02", valid => '1', error => '0'),
        10     => ( data => X"03", valid => '1', error => '0'),
        11     => ( data => X"04", valid => '1', error => '0'),
        12     => ( data => X"05", valid => '1', error => '0'),
        13     => ( data => X"06", valid => '1', error => '0'),
        14     => ( data => X"5A", valid => '1', error => '0'), -- Source Address (5A)
        15     => ( data => X"02", valid => '1', error => '0'),
        16     => ( data => X"03", valid => '1', error => '0'),
        17     => ( data => X"04", valid => '1', error => '0'),
        18     => ( data => X"05", valid => '1', error => '0'),
        19     => ( data => X"06", valid => '1', error => '0'),
        20     => ( data => X"00", valid => '1', error => '0'),
        21     => ( data => X"2E", valid => '1', error => '0'), -- Length/Type = Length = 46
        22     => ( data => X"01", valid => '1', error => '0'),
        23     => ( data => X"02", valid => '1', error => '0'),
        24     => ( data => X"03", valid => '1', error => '0'),
        25     => ( data => X"04", valid => '1', error => '0'),
        26     => ( data => X"05", valid => '1', error => '0'),
        27     => ( data => X"06", valid => '1', error => '0'),
        28     => ( data => X"07", valid => '1', error => '0'),
        29     => ( data => X"08", valid => '1', error => '0'),
        30     => ( data => X"09", valid => '1', error => '0'),
        31     => ( data => X"0A", valid => '1', error => '0'),
        32     => ( data => X"0B", valid => '1', error => '0'),
        33     => ( data => X"0C", valid => '1', error => '0'),
        34     => ( data => X"0D", valid => '1', error => '0'),
        35     => ( data => X"0E", valid => '1', error => '0'),
        36     => ( data => X"0F", valid => '1', error => '0'),
        37     => ( data => X"10", valid => '1', error => '0'),
        38     => ( data => X"11", valid => '1', error => '0'),
        39     => ( data => X"12", valid => '1', error => '0'),
        40     => ( data => X"13", valid => '1', error => '0'),
        41     => ( data => X"14", valid => '1', error => '0'),
        42     => ( data => X"15", valid => '1', error => '0'),
        43     => ( data => X"16", valid => '1', error => '0'),
        44     => ( data => X"17", valid => '1', error => '0'),
        45     => ( data => X"18", valid => '1', error => '0'),
        46     => ( data => X"19", valid => '1', error => '0'),
        47     => ( data => X"1A", valid => '1', error => '0'),
        48     => ( data => X"1B", valid => '1', error => '0'),
        49     => ( data => X"1C", valid => '1', error => '0'),
        50     => ( data => X"1D", valid => '1', error => '0'),
        51     => ( data => X"1E", valid => '1', error => '0'),
        52     => ( data => X"1F", valid => '1', error => '0'),
        53     => ( data => X"20", valid => '1', error => '0'),
        54     => ( data => X"21", valid => '1', error => '0'),
        55     => ( data => X"22", valid => '1', error => '0'),
        56     => ( data => X"23", valid => '1', error => '0'),
        57     => ( data => X"24", valid => '1', error => '0'),
        58     => ( data => X"25", valid => '1', error => '0'),
        59     => ( data => X"26", valid => '1', error => '0'),
        60     => ( data => X"27", valid => '1', error => '0'),
        61     => ( data => X"28", valid => '1', error => '0'),
        62     => ( data => X"29", valid => '1', error => '0'),
        63     => ( data => X"2A", valid => '1', error => '0'),
        64     => ( data => X"2B", valid => '1', error => '0'),
        65     => ( data => X"2C", valid => '1', error => '0'),
        66     => ( data => X"2D", valid => '1', error => '0'),
        67     => ( data => X"2E", valid => '1', error => '0'),
        68     => ( data => X"14", valid => '1', error => '0'), -- FCS field
        69     => ( data => X"19", valid => '1', error => '0'),
        70     => ( data => X"D1", valid => '1', error => '0'),
        71     => ( data => X"DD", valid => '1', error => '0'),
        others => ( data => X"00", valid => '0', error => '0'))
      ),
    1          => (                     -- Frame 1
      columns  => (
        0      => ( data => X"55", valid => '1', error => '0'), -- preamble
        1      => ( data => X"55", valid => '1', error => '0'),
        2      => ( data => X"55", valid => '1', error => '0'),
        3      => ( data => X"55", valid => '1', error => '0'),
        4      => ( data => X"55", valid => '1', error => '0'),
        5      => ( data => X"55", valid => '1', error => '0'),
        6      => ( data => X"55", valid => '1', error => '0'),
        7      => ( data => X"D5", valid => '1', error => '0'), -- SFD
        8      => ( data => X"DA", valid => '1', error => '0'), -- Destination Address (DA)
        9      => ( data => X"02", valid => '1', error => '0'),
        10     => ( data => X"03", valid => '1', error => '0'),
        11     => ( data => X"04", valid => '1', error => '0'),
        12     => ( data => X"05", valid => '1', error => '0'),
        13     => ( data => X"06", valid => '1', error => '0'),
        14     => ( data => X"5A", valid => '1', error => '0'), -- Source Address (5A)
        15     => ( data => X"02", valid => '1', error => '0'),
        16     => ( data => X"03", valid => '1', error => '0'),
        17     => ( data => X"04", valid => '1', error => '0'),
        18     => ( data => X"05", valid => '1', error => '0'),
        19     => ( data => X"06", valid => '1', error => '0'),
        20     => ( data => X"80", valid => '1', error => '0'), -- Length/Type = Type = 8000
        21     => ( data => X"00", valid => '1', error => '0'),
        22     => ( data => X"01", valid => '1', error => '0'),
        23     => ( data => X"02", valid => '1', error => '0'),
        24     => ( data => X"03", valid => '1', error => '0'),
        25     => ( data => X"04", valid => '1', error => '0'),
        26     => ( data => X"05", valid => '1', error => '0'),
        27     => ( data => X"06", valid => '1', error => '0'),
        28     => ( data => X"07", valid => '1', error => '0'),
        29     => ( data => X"08", valid => '1', error => '0'),
        30     => ( data => X"09", valid => '1', error => '0'),
        31     => ( data => X"0A", valid => '1', error => '0'),
        32     => ( data => X"0B", valid => '1', error => '0'),
        33     => ( data => X"0C", valid => '1', error => '0'),
        34     => ( data => X"0D", valid => '1', error => '0'),
        35     => ( data => X"0E", valid => '1', error => '0'),
        36     => ( data => X"0F", valid => '1', error => '0'),
        37     => ( data => X"10", valid => '1', error => '0'),
        38     => ( data => X"11", valid => '1', error => '0'),
        39     => ( data => X"12", valid => '1', error => '0'),
        40     => ( data => X"13", valid => '1', error => '0'),
        41     => ( data => X"14", valid => '1', error => '0'),
        42     => ( data => X"15", valid => '1', error => '0'),
        43     => ( data => X"16", valid => '1', error => '0'),
        44     => ( data => X"17", valid => '1', error => '0'),
        45     => ( data => X"18", valid => '1', error => '0'),
        46     => ( data => X"19", valid => '1', error => '0'),
        47     => ( data => X"1A", valid => '1', error => '0'),
        48     => ( data => X"1B", valid => '1', error => '0'),
        49     => ( data => X"1C", valid => '1', error => '0'),
        50     => ( data => X"1D", valid => '1', error => '0'),
        51     => ( data => X"1E", valid => '1', error => '0'),
        52     => ( data => X"1F", valid => '1', error => '0'),
        53     => ( data => X"20", valid => '1', error => '0'),
        54     => ( data => X"21", valid => '1', error => '0'),
        55     => ( data => X"22", valid => '1', error => '0'),
        56     => ( data => X"23", valid => '1', error => '0'),
        57     => ( data => X"24", valid => '1', error => '0'),
        58     => ( data => X"25", valid => '1', error => '0'),
        59     => ( data => X"26", valid => '1', error => '0'),
        60     => ( data => X"27", valid => '1', error => '0'),
        61     => ( data => X"28", valid => '1', error => '0'),
        62     => ( data => X"29", valid => '1', error => '0'),
        63     => ( data => X"2A", valid => '1', error => '0'),
        64     => ( data => X"2B", valid => '1', error => '0'),
        65     => ( data => X"2C", valid => '1', error => '0'),
        66     => ( data => X"2D", valid => '1', error => '0'),
        67     => ( data => X"2E", valid => '1', error => '0'),
        68     => ( data => X"2F", valid => '1', error => '0'),
        69     => ( data => X"33", valid => '1', error => '0'), -- FCS field
        70     => ( data => X"A9", valid => '1', error => '0'),
        71     => ( data => X"AF", valid => '1', error => '0'),
        72     => ( data => X"1D", valid => '1', error => '0'),
       others  => ( data => X"00", valid => '0', error => '0'))
      ),
    2          => (                     -- Frame 2
     columns   => (
        0      => ( data => X"55", valid => '1', error => '0'), -- preamble
        1      => ( data => X"55", valid => '1', error => '0'),
        2      => ( data => X"55", valid => '1', error => '0'),
        3      => ( data => X"55", valid => '1', error => '0'),
        4      => ( data => X"55", valid => '1', error => '0'),
        5      => ( data => X"55", valid => '1', error => '0'),
        6      => ( data => X"55", valid => '1', error => '0'),
        7      => ( data => X"D5", valid => '1', error => '0'), -- SFD
        8      => ( data => X"DA", valid => '1', error => '0'), -- Destination Address (DA)
        9      => ( data => X"02", valid => '1', error => '0'),
        10     => ( data => X"03", valid => '1', error => '0'),
        11     => ( data => X"04", valid => '1', error => '0'),
        12     => ( data => X"05", valid => '1', error => '0'),
        13     => ( data => X"06", valid => '1', error => '0'),
        14     => ( data => X"5A", valid => '1', error => '0'), -- Source Address (5A)
        15     => ( data => X"02", valid => '1', error => '0'),
        16     => ( data => X"03", valid => '1', error => '0'),
        17     => ( data => X"04", valid => '1', error => '0'),
        18     => ( data => X"05", valid => '1', error => '0'),
        19     => ( data => X"06", valid => '1', error => '0'),
        20     => ( data => X"00", valid => '1', error => '0'),
        21     => ( data => X"2E", valid => '1', error => '0'), -- Length/Type = Length = 46
        22     => ( data => X"01", valid => '1', error => '0'),
        23     => ( data => X"02", valid => '1', error => '0'),
        24     => ( data => X"03", valid => '1', error => '0'),
        25     => ( data => X"04", valid => '1', error => '0'),
        26     => ( data => X"05", valid => '1', error => '0'),
        27     => ( data => X"06", valid => '1', error => '0'),
        28     => ( data => X"07", valid => '1', error => '0'),
        29     => ( data => X"08", valid => '1', error => '0'),
        30     => ( data => X"09", valid => '1', error => '0'),
        31     => ( data => X"0A", valid => '1', error => '0'),
        32     => ( data => X"0B", valid => '1', error => '0'),
        33     => ( data => X"0C", valid => '1', error => '0'),
        34     => ( data => X"0D", valid => '1', error => '0'),
        35     => ( data => X"0E", valid => '1', error => '0'),
        36     => ( data => X"0F", valid => '1', error => '0'),
        37     => ( data => X"10", valid => '1', error => '0'),
        38     => ( data => X"11", valid => '1', error => '0'),
        39     => ( data => X"12", valid => '1', error => '0'),
        40     => ( data => X"13", valid => '1', error => '0'),
        41     => ( data => X"14", valid => '1', error => '0'),
        42     => ( data => X"15", valid => '1', error => '0'),
        43     => ( data => X"16", valid => '1', error => '0'),
        44     => ( data => X"17", valid => '1', error => '0'),
        45     => ( data => X"18", valid => '1', error => '0'),
        46     => ( data => X"19", valid => '1', error => '0'),
        47     => ( data => X"1A", valid => '1', error => '1'), -- Signal an Error
        48     => ( data => X"1B", valid => '1', error => '0'),
        49     => ( data => X"1C", valid => '1', error => '0'),
        50     => ( data => X"1D", valid => '1', error => '0'),
        51     => ( data => X"1E", valid => '1', error => '0'),
        52     => ( data => X"1F", valid => '1', error => '0'),
        53     => ( data => X"20", valid => '1', error => '0'),
        54     => ( data => X"21", valid => '1', error => '0'),
        55     => ( data => X"22", valid => '1', error => '0'),
        56     => ( data => X"23", valid => '1', error => '0'),
        57     => ( data => X"24", valid => '1', error => '0'),
        58     => ( data => X"25", valid => '1', error => '0'),
        59     => ( data => X"26", valid => '1', error => '0'),
        60     => ( data => X"27", valid => '1', error => '0'),
        61     => ( data => X"28", valid => '1', error => '0'),
        62     => ( data => X"29", valid => '1', error => '0'),
        63     => ( data => X"2A", valid => '1', error => '0'),
        64     => ( data => X"2B", valid => '1', error => '0'),
        65     => ( data => X"2C", valid => '1', error => '0'),
        66     => ( data => X"2D", valid => '1', error => '0'),
        67     => ( data => X"2E", valid => '1', error => '0'),
        68     => ( data => X"14", valid => '1', error => '0'), -- FCS field
        69     => ( data => X"19", valid => '1', error => '0'),
        70     => ( data => X"D1", valid => '1', error => '0'),
        71     => ( data => X"DD", valid => '1', error => '0'),
      others   => ( data => X"00", valid => '0', error => '0'))
     ),
   3           => (                     -- Frame 3
     columns   => (
        0      => ( data => X"55", valid => '1', error => '0'), -- Preamble
        1      => ( data => X"55", valid => '1', error => '0'),
        2      => ( data => X"55", valid => '1', error => '0'),
        3      => ( data => X"55", valid => '1', error => '0'),
        4      => ( data => X"55", valid => '1', error => '0'),
        5      => ( data => X"55", valid => '1', error => '0'),
        6      => ( data => X"55", valid => '1', error => '0'),
        7      => ( data => X"D5", valid => '1', error => '0'), -- SFD
        8      => ( data => X"DA", valid => '1', error => '0'), -- Destination Address (DA)
        9      => ( data => X"02", valid => '1', error => '0'),
        10     => ( data => X"03", valid => '1', error => '0'),
        11     => ( data => X"04", valid => '1', error => '0'),
        12     => ( data => X"05", valid => '1', error => '0'),
        13     => ( data => X"06", valid => '1', error => '0'),
        14     => ( data => X"5A", valid => '1', error => '0'), -- Source Address (5A)
        15     => ( data => X"02", valid => '1', error => '0'),
        16     => ( data => X"03", valid => '1', error => '0'),
        17     => ( data => X"04", valid => '1', error => '0'),
        18     => ( data => X"05", valid => '1', error => '0'),
        19     => ( data => X"06", valid => '1', error => '0'),
        20     => ( data => X"00", valid => '1', error => '0'),
        21     => ( data => X"03", valid => '1', error => '0'), -- Length/Type = Length = 03
        22     => ( data => X"01", valid => '1', error => '0'), -- Therefore padding is required
        23     => ( data => X"02", valid => '1', error => '0'),
        24     => ( data => X"03", valid => '1', error => '0'),
        25     => ( data => X"00", valid => '1', error => '0'), -- Padding (uses zero value bytes)
        26     => ( data => X"00", valid => '1', error => '0'),
        27     => ( data => X"00", valid => '1', error => '0'),
        28     => ( data => X"00", valid => '1', error => '0'),
        29     => ( data => X"00", valid => '1', error => '0'),
        30     => ( data => X"00", valid => '1', error => '0'),
        31     => ( data => X"00", valid => '1', error => '0'),
        32     => ( data => X"00", valid => '1', error => '0'),
        33     => ( data => X"00", valid => '1', error => '0'),
        34     => ( data => X"00", valid => '1', error => '0'),
        35     => ( data => X"00", valid => '1', error => '0'),
        36     => ( data => X"00", valid => '1', error => '0'),
        37     => ( data => X"00", valid => '1', error => '0'),
        38     => ( data => X"00", valid => '1', error => '0'),
        39     => ( data => X"00", valid => '1', error => '0'),
        40     => ( data => X"00", valid => '1', error => '0'),
        41     => ( data => X"00", valid => '1', error => '0'),
        42     => ( data => X"00", valid => '1', error => '0'),
        43     => ( data => X"00", valid => '1', error => '0'),
        44     => ( data => X"00", valid => '1', error => '0'),
        45     => ( data => X"00", valid => '1', error => '0'),
        46     => ( data => X"00", valid => '1', error => '0'),
        47     => ( data => X"00", valid => '1', error => '0'),
        48     => ( data => X"00", valid => '1', error => '0'),
        49     => ( data => X"00", valid => '1', error => '0'),
        50     => ( data => X"00", valid => '1', error => '0'),
        51     => ( data => X"00", valid => '1', error => '0'),
        52     => ( data => X"00", valid => '1', error => '0'),
        53     => ( data => X"00", valid => '1', error => '0'),
        54     => ( data => X"00", valid => '1', error => '0'),
        55     => ( data => X"00", valid => '1', error => '0'),
        56     => ( data => X"00", valid => '1', error => '0'),
        57     => ( data => X"00", valid => '1', error => '0'),
        58     => ( data => X"00", valid => '1', error => '0'),
        59     => ( data => X"00", valid => '1', error => '0'),
        60     => ( data => X"00", valid => '1', error => '0'),
        61     => ( data => X"00", valid => '1', error => '0'),
        62     => ( data => X"00", valid => '1', error => '0'),
        63     => ( data => X"00", valid => '1', error => '0'),
        64     => ( data => X"00", valid => '1', error => '0'),
        65     => ( data => X"00", valid => '1', error => '0'),
        66     => ( data => X"00", valid => '1', error => '0'),
        67     => ( data => X"00", valid => '1', error => '0'),
        68     => ( data => X"73", valid => '1', error => '0'), -- FCS field
        69     => ( data => X"00", valid => '1', error => '0'),
        70     => ( data => X"75", valid => '1', error => '0'),
        71     => ( data => X"22", valid => '1', error => '0'),
      others   => ( data => X"00", valid => '0', error => '0'))
     ));


  ------------------------------------------------------------------------------
  -- testbench signals
  ------------------------------------------------------------------------------

  -- signals for the Tx monitor following 8B10B decode
  signal tx_pdata         : std_logic_vector(7 downto 0);
  signal tx_is_k          : std_logic;
  signal stim_tx_clk_1000 : std_logic;
  signal stim_tx_clk_100  : std_logic;
  signal stim_tx_clk_10   : std_logic;
  signal stim_tx_clk      : std_logic;                           -- Transmitter clock (stimulus process).
  signal mon_tx_clk       : std_logic;                           -- Transmitter clock (monitor process).

  -- signals for the Rx stimulus prior to 8B10B encode
  signal rx_pdata         : std_logic_vector(7 downto 0);
  signal rx_is_k          : boolean;
  signal rx_even          : std_logic := '1';                    -- Keep track of the even/odd position
  signal rx_rundisp_pos   : boolean := false;                    -- Indicates +ve running disparity
  signal stim_rx_clk      : std_logic;                           -- Receiver clock (stimulus process).
  signal mon_rx_clk       : std_logic;                           -- Receiver clock (monitor process).
  signal clock_enable     : std_logic;                           -- SGMII mode only: Used to create data at different rates
  signal tx_mon_clock_enable     : std_logic;                           -- SGMII mode only: Used to create data at different rates


  signal gmii_rxd_comp       : std_logic_vector(7 downto 0);

begin  -- behav


  ------------------------------------------------------------------------------
  -- Clock drivers
  ------------------------------------------------------------------------------

  p_stim_rx_clk : process        -- drives Rx stimulus clock at 125 MHz
  begin
      stim_rx_clk <= '0';
      wait for 4 ns;
      stim_rx_clk <= '1';
      wait for 4 ns;
  end process p_stim_rx_clk;

  p_stim_tx_clk_1000 : process        -- drives stim_tx_clk_1000 at 125 MHz
  begin
      stim_tx_clk_1000 <= '0';
      wait for 4 ns;
      stim_tx_clk_1000 <= '1';
      wait for 4 ns;
  end process p_stim_tx_clk_1000;

  p_stim_tx_clk_100 : process         -- drives stim_tx_clk_100 at 12.5 MHz
  begin
      stim_tx_clk_100 <= '0';
        wait for 40 ns;
        stim_tx_clk_100 <= '1';
        wait for 40 ns;
  end process p_stim_tx_clk_100;

  p_stim_tx_clk_10 : process          -- drives stim_tx_clk_100 at 1.25 MHz
  begin
      stim_tx_clk_10 <= '0';
        wait for 400 ns;
        stim_tx_clk_10 <= '1';
        wait for 400 ns;
  end process p_stim_tx_clk_10;


  -- Select between 10Mb/s, 100Mb/s and 1Gb/s Tx clock frequencies
  p_sel_tx_freq : process(speed_is_10_100, speed_is_100, stim_tx_clk_1000, stim_tx_clk_100, stim_tx_clk_10)
  begin
    if speed_is_10_100 = '0' then
      stim_tx_clk <= stim_tx_clk_1000;
    else
      if speed_is_100 = '1' then
        stim_tx_clk <= stim_tx_clk_100;
      else
        stim_tx_clk <= stim_tx_clk_10;
      end if;
    end if;
  end process p_sel_tx_freq;

  gmii_tx_clk <= stim_tx_clk;

  p_gtx_clk : process            -- drives GTX_CLK at 125 MHz
  begin
      gtx_clk <= '0';
      wait for 4 ns;
      gtx_clk <= '1';
      wait for 4 ns;
  end process p_gtx_clk;

  p_pma_rx_clk : process         -- drives pma_rx_clk0 and pma_rx_clk1 at 62.5 MHz
  begin
      pma_rx_clk0 <= '0';
      pma_rx_clk1 <= '1';
      wait until stim_rx_clk'event and stim_rx_clk = '0';
      pma_rx_clk0 <= '1';
      pma_rx_clk1 <= '0';
      wait until stim_rx_clk'event and stim_rx_clk = '0';
  end process p_pma_rx_clk;


  -- monitor clock for the GMII receiver.
  mon_rx_clk <= gmii_rx_clk;



  ------------------------------------------------------------------------------
  -- Tx stimulus process. This process will push frames of data into the
  -- GMII transmitter side of the PCS/PMA core.
  ------------------------------------------------------------------------------
  p_tx_stimulus : process
    variable column_index : natural := 0;  -- Column counter within frame
    variable stats_value  : std_logic_vector(63 downto 0);
  begin

    -- Initialize
    gmii_txd    <= X"FF";
    gmii_tx_en  <= '1';
    gmii_tx_er  <= '1';
    wait for 1 ns;
    gmii_txd    <= X"00";
    gmii_tx_en  <= '0';
    gmii_tx_er  <= '0';

    -- Wait for the configuration process to finish
    wait until configuration_finished;

    -- Transmit four frames through the GMII transmit interface.
    --      -- frame 0 = standard frame
    --      -- frame 1 = type frame
    --      -- frame 2 = frame containing an error
    --      -- frame 3 = standard frame with padding
    assert false
      report "Tx Stimulus " & integer'image(INSTANCE_NUMBER) & ": sending 4 frames ..." & cr
      severity note;

    -- Synchronise to the transmitter clock
    wait until stim_tx_clk'event and stim_tx_clk = '0';

    for frame_index in frame_data'low to frame_data'high loop

      column_index := 0;

      -- loop over columns in frame.
      while to_stdulogic(frame_data(frame_index).columns(column_index).valid) /= '0' loop
        gmii_txd    <= to_stdlogicvector(frame_data(frame_index).columns(column_index).data);
        gmii_tx_en  <= to_stdulogic(frame_data(frame_index).columns(column_index).valid);
        gmii_tx_er  <= to_stdulogic(frame_data(frame_index).columns(column_index).error);
        column_index := column_index + 1;
        wait until stim_tx_clk'event and stim_tx_clk = '0';
      end loop;

      -- Clear the data lines.
      gmii_txd   <= (others => '0');
      gmii_tx_en <= '0';
      gmii_tx_er <= '0';

      for j in 0 to 11 loop                                 -- delay to create Inter Packet Gap.
        wait until stim_tx_clk'event and stim_tx_clk = '0';
      end loop; -- j

    end loop;   -- frame_index
    wait;
  end process p_tx_stimulus;



  ------------------------------------------------------------------------------
  -- The Phy side TBI transmitter output from the core is 8B10B decoded.
  ------------------------------------------------------------------------------

  -- The transmitter monitor clock is provided by the TBI
  mon_tx_clk <= pma_tx_clk;


  p_tx_decode : process
    variable tx_code_group_rev : std_logic_vector(9 downto 0);
    variable decoded_data      : std_logic_vector(7 downto 0);
    variable is_k_var          : boolean;
  begin
    loop
      wait until mon_tx_clk'event and mon_tx_clk = '1';

      -- The bits of tx_code_group must be reversed to match the decode_8b10b function
      for i in 0 to 9 loop
         tx_code_group_rev(i) := tx_code_group(9 - i);
      end loop;

      -- Perform 8B10B decoding of the data stream
      decode_8b10b(
        d10  => tx_code_group_rev,
        q8   => decoded_data,
        is_k => is_k_var);

      -- drive the output signals with the results
      tx_pdata <= decoded_data;

      if is_k_var then
        tx_is_k <= '1';
      else
        tx_is_k <= '0';
      end if;

    end loop;

  end process p_tx_decode;


  ------------------------------------------------------------------------------
  -- Tx Monitor process. This process checks the frames coming out
  -- of the transmitter PHY side interface to make sure that they match
  -- those injected into the transmitter GMII.
  ------------------------------------------------------------------------------
  p_tx_monitor : process
    variable f            : frame_typ;       -- temporary frame variable
    variable column_index : natural   := 0;  -- Column counter

  begin

    -- Compare the transmitted frames to the injected frames
    --      -- frame 0 = standard frame
    --      -- frame 1 = type frame
    --      -- frame 2 = frame containing an error
    --      -- frame 3 = standard frame with padding


    -- then get synced up with the clock
    wait until mon_tx_clk'event and mon_tx_clk = '0';
    -- Wait for the configuration process to finish
    wait until configuration_finished;

    -- loop over all the frames in the stimulus vector
    for frame_index in frame_data'low to frame_data'high loop
      column_index := 0;

      -- Detect the Start of Frame
      while tx_pdata /= X"FB" loop -- /K27.7/ character
        wait until mon_tx_clk'event and mon_tx_clk = '0';
      end loop;

      -- Move past the Start of Frame code to the 1st byte of preamble
      wait until mon_tx_clk'event and mon_tx_clk = '0' and tx_mon_clock_enable = '1';

      -- wait until the SFD code is detected.
      -- NOTE: It is neccessary to resynchronise on the SFD as the preamble field
      --       may have shrunk.
      while tx_pdata /= X"D5" loop
          assert (tx_pdata = to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)))
          report "Tx Monitor " & integer'image(INSTANCE_NUMBER) & ": data incorrect during the preamble of frame" & integer'image(frame_index) & cr
          severity error;

        -- wait for next column of data
        column_index := column_index + 1;
        wait until mon_tx_clk'event and mon_tx_clk = '0' and tx_mon_clock_enable = '1';
      end loop;

      -- tx_pdata should now hold the SFD.  We need to move to the SFD of the injected frame.
      while to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)) /= X"D5" loop
        column_index := column_index + 1;
      end loop;

      -- Start comparing transmitted frame data to the injected frame data
      assert false
        report "Tx Monitor " & integer'image(INSTANCE_NUMBER) & ": Comparing transmitted frame " & integer'image(frame_index) &" with injected frame " & integer'image(frame_index) & cr
        severity note;

      -- frame has started, loop over columns of frame until the frame termination is detected
      while tx_pdata /= X"FD" or tx_is_k /= '1' loop -- /K29.7/ character

        if tx_pdata /= X"FE" and tx_is_k /= '1' then            -- Do not check the data if an error code has been inserted (/K30.7 character).
          if tx_mon_clock_enable = '1' then
            assert (tx_pdata = to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)))
              report "Tx frame data: " & integer'image(to_integer(unsigned(tx_pdata))) & ", Tx record data: " & integer'image(to_integer(unsigned(to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0))))) & cr & "Tx Monitor: data incorrect during frame" & integer'image(frame_index) & cr
              severity error;
          end if;
        end if;

        -- wait for next column of data
        if tx_mon_clock_enable = '1' then
          column_index := column_index + 1;
        end if;
        wait until mon_tx_clk'event and mon_tx_clk = '0';
      end loop;
    end loop;  -- frame_index

    wait for 200 ns;
    tx_monitor_finished <= true;

  end process p_tx_monitor;



  ------------------------------------------------------------------------------
  -- Rx stimulus process. This process will create frames of data to be
  -- pushed into the receiver PHY side of the PCS/PMA core.
  ------------------------------------------------------------------------------

  -- Set the expected data rate: sample the data on every clock at
  -- 1Gbps, every 10 clocks at 100Mbps, every 100 clocks at 10Mbps
  rx_sample_gen: process (stim_rx_clk)
    variable sample_count: integer range 0 to 99 := 0;
  begin
    if stim_rx_clk'event and stim_rx_clk = '1' then
      if speed_is_10_100 = '0' then
        sample_count   := 0;
        clock_enable <= '1';                                    -- sample on every clock
      else
        if (speed_is_100 = '1' and  sample_count = 9) or    -- sample every 10 clocks
           (speed_is_100 = '0' and  sample_count = 99) then -- sample every 100 clocks
          sample_count   := 0;
          clock_enable <= '1';
        else
          if (sample_count = 99) then
            sample_count := 0;
          else
            sample_count := sample_count + 1;
          end if;
          clock_enable <= '0';
        end if;
      end if;
      if speed_is_10_100 = '0' then
        tx_mon_clock_enable <= '1';                                    -- sample on every clock
      else
        if (speed_is_100 = '1' and  sample_count = 9) or    -- sample every 10 clocks
           (speed_is_100 = '0' and  sample_count = 99) then -- sample every 100 clocks
          tx_mon_clock_enable <= '1';
        else
          tx_mon_clock_enable <= '0';
        end if;
      end if;

    end if;
  end process rx_sample_gen;


  p_rx_stimulus : process
    variable column_index : natural := 0;  -- Column counter within frame

    -- A procedure to create an Idle /I1/ code group
    procedure send_I1 is
    begin
      rx_pdata  <= X"BC";  -- /K28.5/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
      rx_pdata  <= X"C5";  -- /D5.6/
      rx_is_k   <= false;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
    end send_I1;

    -- A procedure to create an Idle /I2/ code group
    procedure send_I2 is
    begin
      rx_pdata  <= X"BC";  -- /K28.5/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
      rx_pdata  <= X"50";  -- /D16.2/
      rx_is_k   <= false;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
    end send_I2;

    -- A procedure to create a Start of Packet /S/ code group
    procedure send_S is
    begin
      rx_pdata  <= X"FB";  -- /K27.7/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
    end send_S;

    -- A procedure to create a Terminate /T/ code group
    procedure send_T is
    begin
      rx_pdata  <= X"FD";  -- /K29.7/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
    end send_T;

    -- A procedure to create a Carrier Extend /R/ code group
    procedure send_R is
    begin
      rx_pdata  <= X"F7";  -- /K23.7/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1';
    end send_R;

    -- A procedure to create an Error Propogation /V/ code group
    procedure send_V is
    begin
      rx_pdata  <= X"FE";  -- /K30.7/
      rx_is_k   <= true;
      wait until stim_rx_clk'event and stim_rx_clk = '1' and clock_enable = '1';
    end send_V;


  begin

    -- Wait for the Management MDIO transaction to finish.
    while not configuration_finished loop
      send_I2;
    end loop;

    -- Inject four frames into the receiver PHY interface
    --      -- frame 0 = standard frame
    --      -- frame 1 = type frame
    --      -- frame 2 = frame containing an error
    --      -- frame 3 = standard frame with padding
    assert false
      report "Rx Stimulus " & integer'image(INSTANCE_NUMBER) & ": sending 4 frames ... " & cr
      severity note;

    for frame_index in frame_data'low to frame_data'high loop

      ------------------------------------
      -- Send a Start of Packet code group
      ------------------------------------
      send_S;

      ------------------------------------
      -- Send frame data
      ------------------------------------
      column_index := 1;

      -- loop over columns in frame
      while to_stdulogic(frame_data(frame_index).columns(column_index).valid) /= '0' loop
        if to_stdulogic(frame_data(frame_index).columns(column_index).error) = '1' then
          send_V; -- insert an error propogation code group
        else
          rx_pdata    <= to_stdlogicvector(frame_data(frame_index).columns(column_index).data);
          rx_is_k     <= false;
          wait until stim_rx_clk'event and stim_rx_clk = '1' and clock_enable = '1';
        end if;
        column_index := column_index + 1;
      end loop;

      ------------------------------------
      -- Send a frame termination sequence
      ------------------------------------
      send_T;    -- Terminate code group
      send_R;    -- Carrier Extend code group

     -- An extra Carrier Extend code group should be sent to end the frame
     -- on an even boundary.
      if rx_even = '1' then
        send_R;  -- Carrier Extend code group
      end if;

      ------------------------------------
      -- Send an Inter Packet Gap.
      ------------------------------------
     -- The initial Idle following a frame should be chosen to ensure
     -- that the running disparity is returned to -ve.
      if rx_rundisp_pos then
        send_I1;  -- /I1/ will flip the running disparity
      else
        send_I2;  -- /I2/ will maintain the running disparity
      end if;

      -- The remainder of the IPG is made up of /I2/ 's.
      -- NOTE: the number 4 in the following calculations is made up
      --      from 2 bytes of the termination sequence and 2 bytes from
      --      the initial Idle.
      if speed_is_10_100 = '0' then
        for j in 0 to 3 loop       -- 4 /I2/'s = 8 clock periods (12 - 4)
          send_I2;
        end loop; -- j
      else
        if speed_is_100 = '1' then -- 58 /I2/'s = 116 clock periods (120 - 4)
          for j in 0 to 57 loop
            send_I2;
          end loop; -- j
        else
          for j in 0 to 597 loop   -- 598 /I2/'s = 1196 clock periods (1200 - 4)
            send_I2;
          end loop; -- j
        end if;
      end if;

    end loop;   -- frame_index

    -- After the completion of the simulus, send Idles continuously
    loop
      send_I2;
    end loop;

  end process p_rx_stimulus;



  ------------------------------------------------------------------------------
  -- A process to keep track of the even/odd code group position for the
  -- injected receiver code groups.
  ------------------------------------------------------------------------------
  p_rx_even_odd: process
  begin
    wait until stim_rx_clk'event and stim_rx_clk = '1';
    rx_even <= not rx_even;
  end process p_rx_even_odd;


  ------------------------------------------------------------------------------
  -- Data from the Rx Stimulus is 8B10B encoded so that it can be
  -- injected into the TBI receiver port.
  ------------------------------------------------------------------------------
  p_rx_encode : process
    variable encoded_data     : std_logic_vector(9 downto 0) := (others => '0');
    variable encoded_data_rev : std_logic_vector(9 downto 0) := (others => '0');
    variable rundisp          : boolean;
  begin

    -- Drive with initial value
    rx_code_group  <= "0000000000";

    -- Get synced up with the Rx clock
    wait until stim_rx_clk'event and stim_rx_clk = '1';

    loop
    -- Perform 8B10B encoding of the data stream
       encode_8b10b(
         d8                => rx_pdata,
         is_k              => rx_is_k,
         disparity_pos_in  => rundisp,
         q10               => encoded_data,
         disparity_pos_out => rundisp);

       -- The bits of encoded_data must be reversed to match the encode_8b10b function
       for i in 0 to 9 loop
          encoded_data_rev(i) := encoded_data(9 - i);
       end loop;

       -- drive the output signals with the results
       rx_rundisp_pos <= rundisp;
       rx_code_group  <= encoded_data_rev;

       wait until stim_rx_clk'event and stim_rx_clk = '1';
    end loop;

  end process p_rx_encode;



  ------------------------------------------------------------------------------
  -- Rx monitor process. This process checks the data coming out of the
  -- receiver GMII to make sure that it matches that injected into the
  -- PHY.
  ------------------------------------------------------------------------------
  gmii_rxd_comp <= gmii_rxd;

  p_rx_monitor : process
    variable f            : frame_typ;       -- temporary frame variable
    variable column_index : natural   := 0;  -- Column counter

  begin

    -- Compare the received frames to the injected frames
    --      -- frame 0 = standard frame
    --      -- frame 1 = type frame
    --      -- frame 2 = frame containing an error
    --      -- frame 3 = standard frame with padding

    wait for 1 us;

    -- then get synced up with the rx clock
    if gmii_rx_dv /= '0' then
       wait until gmii_rx_dv = '0';
    end if;
    wait until mon_rx_clk'event and mon_rx_clk = '1';

    -- loop over all the frames in the stimulus vector
    for frame_index in frame_data'low to frame_data'high loop
      column_index := 0;

      -- wait for the first real column of data to come out of Rx GMII
      while gmii_rx_dv = '0' loop
    wait until mon_rx_clk'event and mon_rx_clk = '1';
      end loop;


      -- wait until the SFD code is detected on gmii_rxd(7 downto 0).
      -- NOTE: It is neccessary to resynchronise on the SFD as the preamble field
      --       may have shrunk.
      while gmii_rxd_comp /= X"D5" loop
        assert (gmii_rx_dv = to_stdUlogic(frame_data(frame_index).columns(column_index).valid))
          report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rx_dv incorrect during the preamble of frame " & integer'image(frame_index) & cr
          severity error;

        assert (gmii_rx_er = to_stdUlogic(frame_data(frame_index).columns(column_index).error))
          report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rx_er incorrect during the preamble of frame " & integer'image(frame_index) & cr
          severity error;

        assert (gmii_rxd_comp(7 downto 0) =
                to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)))
          report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rxd incorrect during the preamble of frame " & integer'image(frame_index) & cr
          severity error;

        -- wait for next column of data
        column_index := column_index + 1;
        wait until mon_rx_clk'event and mon_rx_clk = '1';

      end loop;


      -- gmii_rxd should now hold the SFD.  We need to move to the SFD of the injected frame.
      while to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)) /= X"D5" loop
        column_index := column_index + 1;
      end loop;

      -- Start comparing received data to injected data
      assert false
        report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": Comparing received frame " & integer'image(frame_index) &" with injected frame " & integer'image(frame_index) & cr
        severity note;

      -- frame has started, loop over columns of frame
      while gmii_rx_dv /= to_stdUlogic('0') loop
          assert (gmii_rx_dv = to_stdUlogic(frame_data(frame_index).columns(column_index).valid))
            report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rx_dv incorrect during frame " & integer'image(frame_index) & cr
            severity error;

          assert (gmii_rx_er = to_stdUlogic(frame_data(frame_index).columns(column_index).error))
            report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rx_er incorrect during frame " & integer'image(frame_index) & cr
            severity error;

          if gmii_rx_er = '0' then            -- Do not check the data if an error code has been inserted.
            assert (gmii_rxd_comp(7 downto 0) =
                    to_stdlogicvector(frame_data(frame_index).columns(column_index).data(7 downto 0)))
              report "Rx Monitor " & integer'image(INSTANCE_NUMBER) & ": gmii_rxd incorrect during frame " & integer'image(frame_index) & cr
              severity error;
          end if;

        -- wait for next column of data
        column_index := column_index + 1;
        wait until mon_rx_clk'event and mon_rx_clk = '1';
      end loop;  -- while data valid
    end loop;  -- frame_index

    wait for 200 ns;
    rx_monitor_finished <= true;

  end process p_rx_monitor;



end behav;

